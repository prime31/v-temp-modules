module yoga

#flag -I @VMOD/prime31/yoga/thirdparty
#flag darwin @VMOD/prime31/yoga/thirdparty/libyogacore.a
#flag darwin -lc++

#flag linux @VMOD/prime31/yoga/thirdparty/libyogacore.a
#flag linux -lstdc++

#include "Yoga.h"
