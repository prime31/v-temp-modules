module mixer
