module fmod
import prime31.fmod.core

struct Dsp {
pub:
	dsp &FMOD_DSP
}