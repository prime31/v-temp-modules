module fmod

struct Dsp {
pub:
	dsp &FMOD_DSP
}