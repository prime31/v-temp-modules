module gl3w

