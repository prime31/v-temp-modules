module truetype

#flag -I @VMOD/prime31/stb/truetype/thirdparty

#define STB_RECT_PACK_IMPLEMENTATION
#include "stb_rect_pack.h"

#define STB_TRUETYPE_IMPLEMENTATION 
#include "stb_truetype.h"

