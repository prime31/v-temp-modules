module sdl2_image