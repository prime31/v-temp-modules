module physfs

