module fmod

pub struct SoundGroup {
pub:
	group &FMOD_SOUNDGROUP
}