module via

struct Audio {
	
}

fn create_audio(config ViaConfig) &Audio {
	return &Audio{}
}