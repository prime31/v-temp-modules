module fmod
import prime31.fmod.core

pub struct SoundGroup {
pub:
	group &FMOD_SOUNDGROUP
}