module core

struct Dsp {
pub:
	dsp &FMOD_DSP
}