module sokol
import prime31.sokol.c


