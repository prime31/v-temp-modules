module ttf

