module via

struct Timer {
	
}

fn create_timer(config ViaConfig) &Timer {
	return &Timer{}
}