module gl3w

fn C.gl3wInit()