module sdl2_mixer
