module gl3w

pub fn initialize() {
	C.gl3wInit()
}