module image