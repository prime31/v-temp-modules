module via

struct FileSystem {
	
}

fn create_filesystem(config ViaConfig) &FileSystem {
	return &FileSystem{}
}