module via

struct Graphics {
	
}

fn create_graphics(config ViaConfig) &Graphics {
	return &Graphics{}
}