module via

struct Window {
	
}

fn create_window(config ViaConfig) &Window {
	return &Window{}
}