module image
