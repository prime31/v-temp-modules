module sdl2_ttf

