module physfs


#flag -I @VMOD/prime31/physfs/physfs_hg/src
#flag darwin -framework IOKit -framework Foundation
#flag darwin @VMOD/prime31/physfs/physfs_hg/build/libphysfs.a

#include "physfs.h"
