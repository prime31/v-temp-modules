module physfs_impl


